`timescale 1ps/1ps
`include "command_FSM_if.vh"

module command_FSM (
    input logic CLK,
    input logic nRST,
    command_FSM_if.dut mycmd
);
    import dram_pkg::*;
    localparam logic [1:0] IDLE_R = 2'b00;
    localparam logic [1:0] HIT = 2'b01;
    localparam logic [1:0] MISS = 2'b10;
    localparam logic [1:0] CONFLICT = 2'b11;
    logic nram_wait;

    always_ff @(posedge CLK, negedge nRST) begin
        if (!nRST) begin
            mycmd.cmd_state <= POWER_UP;
        end else begin
            mycmd.cmd_state <= mycmd.ncmd_state;
        end
    end

    always_ff @(posedge CLK, negedge nRST) begin
        if (!nRST) begin
            mycmd.ram_wait <= 1;
        end else begin
            mycmd.ram_wait <= nram_wait;
        end
    end

    always_comb begin
        mycmd.ncmd_state = mycmd.cmd_state;
        mycmd.row_resolve = 1'b0;
        mycmd.init_req = 0;
        nram_wait = 1;
        casez (mycmd.cmd_state)

            POWER_UP: begin
                mycmd.init_req = 1;
                if (mycmd.init_done) mycmd.ncmd_state = IDLE;
            end

            REFRESH: begin
                mycmd.ncmd_state = REFRESHING;
                
            end

            REFRESHING: begin
                if (mycmd.tREF_done) begin
                    mycmd.ncmd_state = IDLE;     
                end
            end

            IDLE: begin
                if (mycmd.rf_req) begin
                    // mycmd.ncmd_state = (mycmd.all_row_closed) ? REFRESH : PRECHARGE;
                    mycmd.ncmd_state = PRECHARGE_RE;
                end
                else if (mycmd.dWEN || mycmd.dREN) begin
                    if (mycmd.row_stat == HIT) mycmd.ncmd_state = mycmd.dWEN ? WRITE : READ;
                    else if(mycmd.row_stat == CONFLICT) mycmd.ncmd_state = PRECHARGE;
                    else if (mycmd.row_stat == MISS) mycmd.ncmd_state = ACTIVATE;
                end
            end

            ACTIVATE: begin
                // if (mycmd.rf_req) begin mycmd.ncmd_state = (mycmd.all_row_closed) ? REFRESH : PRECHARGE; end
                if (mycmd.rf_req) begin mycmd.ncmd_state = PRECHARGE_RE; end
                else begin mycmd.ncmd_state = ACTIVATING; end
            end

            ACTIVATING: begin
                if (mycmd.tACT_done) begin
                    mycmd.ncmd_state = mycmd.rf_req ? PRECHARGE_RE : mycmd.dWEN ? WRITE : READ;
                end
            end

            WRITE: begin mycmd.ncmd_state = mycmd.rf_req ? PRECHARGE_RE : WRITING; end
            READ : begin mycmd.ncmd_state = mycmd.rf_req ? PRECHARGE_RE : READING; end
            
            WRITING: begin
                if (mycmd.tWR_done) begin
                    nram_wait = 1'b0;
                    if (mycmd.rf_req) begin mycmd.ncmd_state = PRECHARGE_RE; end
                    //TODO Discuss this with Dhruv
                    // else if (mycmd.dWEN || mycmd.dREN) begin
                    //     if (mycmd.row_stat == HIT) mycmd.ncmd_state = mycmd.dWEN ? WRITE : READ;
                    //     else if(mycmd.row_stat == CONFLICT) mycmd.ncmd_state = PRECHARGE;
                    //     else if (mycmd.row_stat == MISS) mycmd.ncmd_state = ACTIVATE;
                    // end 
                    else begin
                        mycmd.ncmd_state = IDLE;
                    end 
                end
            end

            READING: begin
                if (mycmd.tRD_done) begin
                    nram_wait = 1'b0;
                    if (mycmd.rf_req) begin mycmd.ncmd_state = PRECHARGE_RE; end
                    //TODO Discuss this with Dhruv
                    // else if [(mycmd.dWEN || mycmd.dREN) begin
                    //     if (mycmd.row_stat == HIT) mycmd.ncmd_state = mycmd.dWEN ? WRITE : READ;
                    //     else if(mycmd.row_stat == CONFLICT) mycmd.ncmd_state = PRECHARGE;
                    //     else if (mycmd.row_stat == MISS) mycmd.ncmd_state = ACTIVATE;
                    // end
                    else begin
                        mycmd.ncmd_state = IDLE;
                    end 
                end 
            end

            PRECHARGE: begin
                mycmd.ncmd_state = PRECHARGING;
            end

            PRECHARGING: begin
                if (mycmd.tPRE_done) begin
                    mycmd.row_resolve = 1'b1;
                    if (mycmd.rf_req) begin
                        mycmd.ncmd_state = PRECHARGE_RE;    
                    end else begin
                        mycmd.ncmd_state = IDLE;
                    end
                end
            end

            PRECHARGE_RE: begin
                mycmd.ncmd_state = PRECHARGING_RE;
            end

            PRECHARGING_RE: begin
                if (mycmd.tPRE_done) begin
                    mycmd.ncmd_state = REFRESH;
                end
            end
        endcase
    end

endmodule
