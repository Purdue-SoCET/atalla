`include "sqrt_types.vh"
`include "sqrt_fp16_if.sv"

module sqrt_bf16 (
    input logic         CLK,
    input logic         nRST,
    sqrt_if.srif        srif
)

    


endmodule