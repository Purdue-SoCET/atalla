80'b00000000000000000000000000000000000000000000000000000000000000000000000000000000,
80'b11111111111111110101010101010101000100010001000100000001000000010000000000000001,
80'b00000000000000001111111111111111001100110011001100000011000000110000000000000011,
80'b11111111111111111010101010101010011101110111011100000111000001110000000000000111,
80'b00000000000000000000000000000000111111111111111100001111000011110000000000001111,
80'b11111111111111110101010101010101111011101110111000011111000111110000000000011111,
80'b00000000000000001111111111111111110011001100110000111111001111110000000000111111,
80'b11111111111111111010101010101010100010001000100001111111011111110000000001111111,
80'b00000000000000000000000000000000000000000000000011111111111111110000000011111111,
80'b11111111111111110101010101010101000100010001000111111110111111100000000111111111,
80'b00000000000000001111111111111111001100110011001111111100111111000000001111111111,
80'b11111111111111111010101010101010011101110111011111111000111110000000011111111111,
80'b00000000000000000000000000000000111111111111111111110000111100000000111111111111,
80'b11111111111111110101010101010101111011101110111011100000111000000001111111111111,
80'b00000000000000001111111111111111110011001100110011000000110000000011111111111111,
80'b11111111111111111010101010101010100010001000100010000000100000000111111111111111,
80'b00000000000000000000000000000000000000000000000000000000000000001111111111111111,
80'b11111111111111110101010101010101000100010001000100000001000000011111111111111110,
80'b00000000000000001111111111111111001100110011001100000011000000111111111111111100,
80'b11111111111111111010101010101010011101110111011100000111000001111111111111111000,
80'b00000000000000000000000000000000111111111111111100001111000011111111111111110000,
80'b11111111111111110101010101010101111011101110111000011111000111111111111111100000,
80'b00000000000000001111111111111111110011001100110000111111001111111111111111000000,
80'b11111111111111111010101010101010100010001000100001111111011111111111111110000000,
80'b00000000000000000000000000000000000000000000000011111111111111111111111100000000,
80'b11111111111111110101010101010101000100010001000111111110111111101111111000000000,
80'b00000000000000001111111111111111001100110011001111111100111111001111110000000000,
80'b11111111111111111010101010101010011101110111011111111000111110001111100000000000,
80'b00000000000000000000000000000000111111111111111111110000111100001111000000000000,
80'b11111111111111110101010101010101111011101110111011100000111000001110000000000000,
80'b00000000000000001111111111111111110011001100110011000000110000001100000000000000,
80'b11111111111111111010101010101010100010001000100010000000100000001000000000000000