`ifndef DRAM_PKG_VH
`define DRAM_PKG_VH

package dram_pkg;

    // WORD SIZE
    parameter WORD_W            = 32;

    // CONFIGS
    parameter CONFIG_BITS = 2;
    
    // ADDRESS PARAMETERS
    parameter RANK_BITS         = 1;
    parameter BANK_GROUP_BITS   = 2;
    parameter BANK_BITS         = 2;
    parameter ROW_BITS          = 15;
    parameter COLUMN_BITS       = 10;
    parameter OFFSET_BITS       = 2;
    parameter IGNORE_BITS       = 1;
    parameter ADDR_BITS         = 14;

    // TIMING PARAMETERS
    parameter tRCD = 10;
    parameter tAL = 0;
    parameter tCL = 10;
    parameter tBURST = 4;
    parameter tCWL = 10;
    parameter tREFI = 250;
    parameter tRP = 10;
    parameter tRFC = 172;
    parameter tRAS = 45;
    parameter tRC = tRAS + tRP;
    parameter tRL = tAL + tCL;        // Read Latency
    parameter tWL = tAL + tCWL;       // Write Latency
    parameter MAX_tREFRESH_LIMIT = 9 * tREFI;
    parameter tWR = 13;
    parameter tWTR = 5;

    //INITIALIZE TIMING PARAMETERS
    parameter tRESET        = 80;
    parameter tPWUP         = 80;
    parameter tRESETCKE     = 80;
    parameter tPDc          = 3;
    parameter tXPR          = 217;
    parameter tDLLKc        = 597;
    parameter tZQinitc      = 1024;
    parameter tMOD          = 25;

    // word_t
    typedef logic [WORD_W-1:0] word_t;

    // configs_t - x4, x8, x16
    typedef enum logic [CONFIG_BITS-1:0] {
        x4  = 2'b00,
        x8  = 2'b01,
        x16 = 2'b10
    } configs_t;

    // DRAM init/command states
    typedef enum logic [4:0] {
        POWER_UP,
        PRE_RESET,
        RESET,
        NOP,
        LOAD_MODE_DLL,
        LOAD_BG0_REG3,
        LOAD_BG1_REG6,
        LOAD_BG1_REG5,
        LOAD_BG1_REG4,
        LOAD_BG0_REG2,
        LOAD_BG0_REG1,
        LOAD_BG0_REG0,
        ZQ_CL,
        IDLE,
        ACTIVATE,
        ACTIVATING,
        WRITE,
        WRITING,
        PRECHARGE,
        PRECHARGING,
        PRECHARGING_ALL,
        READ,
        READING,
        REFRESH,
        REFRESHING
    } dram_state_t; 

    // {cs, act, ras, cas, we}
    typedef enum logic [4:0] {
        POWER_UP_PRG  = 5'b01111,
        LOAD_MODE_CMD = 5'b01000,
        REFRESH_CMD   = 5'b01001,
        PRECHARGE_CMD = 5'b01010,
        ACTIVATE_CMD  = 5'b00xxx,
        WRITE_CMD     = 5'b01100,
        READ_CMD      = 5'b01101,
        ZQ_CMD        = 5'b01110,
        DESEL_CMD     = 5'b11000
    } cmd_t;

    // DRAM CONFIGURATIONS
    parameter BURST_LENGTH  = 8;
    parameter CONFIGURED_DQ_BITS     = 16;
    parameter CONFIGURED_DQS_BITS     = 16;
    parameter CONFIGURED_DM_BITS     = 16;
    parameter CONFIGURED_RANKS = 1;
    parameter DM_BITS       = 16;

endpackage

`endif // DRAM_PKG_VH