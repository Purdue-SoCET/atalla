
`timescale 1ns/1ps

module wallacetree_11b_mini #(parameter NUM_BITS = 11) (input logic [10:0] a, b, output logic [12:0] result, output logic overflow, round_loss, output logic [21:0] debug_output);

    // I have no idea if this works for NUM_BITS other than 11. ceil(11/2)is 6, but since indices are 0 indexed in Verilog, I am using floor(11/2) which is 5 so perfect for [5:0]

    logic [NUM_BITS+1:0] extended_multiplier;
    logic [NUM_BITS/2:0][2:0] booth_multipliers;

    genvar z, x, c, v;

    // Generate multiplier chunks
    assign extended_multiplier = {1'b0, b, 1'b0};       // Put a 0 at the MSB and LSB of multiplier (b)
    generate
        for(z = 0; z <= NUM_BITS / 2; z++)
        begin
            assign booth_multipliers[z] = extended_multiplier[ (z*2)+2 : (z*2) ];
        end
    endgenerate

    // Generate partial products
    // Logic from here: https://ieeexplore.ieee.org/document/9121226
    // logic written with GPT edits
    logic signed [NUM_BITS/2 : 0][NUM_BITS+1:0] pprod;      // each partial product should be 2 bits longer than the input, to accommodate an input left-shifted by 1 and a sign bit.
    generate
        for(x = 0; x <= NUM_BITS/2; x++)
        begin
            // logic: if the booth encoded multiplier chunk is negative (MSB is 1), set the partial product to -(value << [the magnitude of the multiplier chunk]). Else, just set it to (value << [the magnitude of the multiplier chunk]). Negation is done with 2's complement: invert bits and add 1.
            always_comb begin
                casez(booth_multipliers[x])
                    3'b000, 3'b111: pprod[x] = '0;

                    3'b001, 3'b010: pprod[x] = {2'b00, a};
                    3'b011: pprod[x] = {1'b0, a} << 1;

                    3'b101, 3'b110: pprod[x] = (~{2'b00, a}) + 1;
                    3'b100: pprod[x] = ~({1'b0, a, 1'b0}) + 1;
                endcase
            end
        end
    endgenerate

    // 11 by 6 wallace tree. we only have 6 partial products.

    // layer 1: 4:2 compressors compressing partial products 0 through 3
    logic [18:0] level1_sums;
    logic [14:0] level1_carries;
    logic [9:0] level1_internal_carries;

    // sum[1:0] assigned directly from pp0
    assign level1_sums[1:0] = pprod[0][1:0];

    // sum[3:2] halfadders
    ha ha_l1_b2(.a(pprod[0][2]), .b(pprod[1][0]), .s(level1_sums[2]), .cout(level1_carries[0]));
    ha ha_l1_b3(.a(pprod[0][3]), .b(pprod[1][1]), .s(level1_sums[3]), .cout(level1_carries[1]));

    // sum[5:4] full adders 
    fa fa_l1_b4(.a(pprod[0][4]), .b(pprod[1][2]), .cin(pprod[2][0]), .s(level1_sums[4]), .cout(level1_carries[2]));
    fa fa_l1_b5(.a(pprod[0][5]), .b(pprod[1][3]), .cin(pprod[2][1]), .s(level1_sums[5]), .cout(level1_carries[3]));

    // sum[12:6] 4:2 compressors
    assign level1_internal_carries[0] = 1'b0;   // first 4:2 compressor has no carry in
    generate
        for(c = 6; c <= 12; c++)
        begin
            compress_4to2 c42_l1(.x1(pprod[0][c]), .x2(pprod[1][c-2]), .x3(pprod[2][c-4]), .x4(pprod[3][c-6]), .cin(level1_internal_carries[c-6]), .sum(level1_sums[c]), .carry(level1_carries[c-2]), .cout(level1_internal_carries[c-5]));
        end
    endgenerate

    //sum[14:13] 4:2 compressors with x1=0
    compress_4to2 c42_l1_b13(.x1(1'b0), .x2(pprod[1][11]), .x3(pprod[2][9]), .x4(pprod[3][7]), .cin(level1_internal_carries[7]), .sum(level1_sums[13]), .carry(level1_carries[11]), .cout(level1_internal_carries[8]));
    compress_4to2 c42_l1_b14(.x1(1'b0), .x2(pprod[1][12]), .x3(pprod[2][10]), .x4(pprod[3][8]), .cin(level1_internal_carries[8]), .sum(level1_sums[14]), .carry(level1_carries[12]), .cout(level1_internal_carries[9]));

    //sum[15] full adder. must be a fa not an ha to deal with the carry generated by the 4:2 compressor
    fa fa_l1_b15(.a(level1_internal_carries[9]), .b(pprod[2][11]), .cin(pprod[3][9]), .s(level1_sums[15]), .cout(level1_carries[13]));

    //sum[16] half adder
    ha ha_l1_b16(.a(pprod[2][12]), .b(pprod[3][10]), .s(level1_sums[16]), .cout(level1_carries[14]));

    //sum[18:17] assigned directly from pp3
    assign level1_sums[18:17] = pprod[3][12:11];



    // layer 2: more 4:2 compressors compressing the 2 lines from level1 and the remaining 2 partial products
    logic [22:0] level2_sums;
    logic [17:0] level2_carries;
    logic [9:0] level2_internal_carries;

    // sum[2:0] assigned directly from previous layer
    assign level2_sums[2:0] = level1_sums[2:0];

    // sum[7:3] halfadders
    ha ha_l2_b3(.a(level1_sums[3]), .b(level1_carries[0]), .s(level2_sums[3]), .cout(level2_carries[0]));
    ha ha_l2_b4(.a(level1_sums[4]), .b(level1_carries[1]), .s(level2_sums[4]), .cout(level2_carries[1]));
    ha ha_l2_b5(.a(level1_sums[5]), .b(level1_carries[2]), .s(level2_sums[5]), .cout(level2_carries[2]));
    ha ha_l2_b6(.a(level1_sums[6]), .b(level1_carries[3]), .s(level2_sums[6]), .cout(level2_carries[3]));
    ha ha_l2_b7(.a(level1_sums[7]), .b(level1_carries[4]), .s(level2_sums[7]), .cout(level2_carries[4]));

    // sum[9:8] fulladders
    fa fa_l2_b8(.a(level1_sums[8]), .b(level1_carries[5]), .cin(pprod[4][0]), .s(level2_sums[8]), .cout(level2_carries[5]));
    fa fa_l2_b9(.a(level1_sums[9]), .b(level1_carries[6]), .cin(pprod[4][1]), .s(level2_sums[9]), .cout(level2_carries[6]));

    // sum[17:10] 4:2 compressors
    assign level2_internal_carries[0] = 1'b0;
    generate
        for(v = 10; v <= 17; v++)
        begin
            compress_4to2 c42_l2(.x1(pprod[4][v-8]), .x2(pprod[5][v-10]), .x3(level1_sums[v]), .x4(level1_carries[v-3]), .cin(level2_internal_carries[v-10]), .sum(level2_sums[v]), .carry(level2_carries[v-3]), .cout(level2_internal_carries[v-9]));
        end
    endgenerate

    // sum[18] 4:2 compressor with x4=0
    compress_4to2 c42_l2_b18(.x1(pprod[4][10]), .x2(pprod[5][8]), .x3(level1_sums[18]), .x4(1'b0), .cin(level2_internal_carries[8]), .sum(level2_sums[18]), .carry(level2_carries[15]), .cout(level2_internal_carries[9]));

    // sum[19] full adder
    fa fa_l2_b19(.a(level2_internal_carries[9]), .b(pprod[4][11]), .cin(pprod[5][9]), .s(level2_sums[19]), .cout(level2_carries[16]));
    
    // sum[20] half adder
    ha ha_l2_b20(.a(pprod[4][12]), .b(pprod[5][10]), .s(level2_sums[20]), .cout(level2_carries[17]));

    // sum[22:21] assigned directly from pp5
    assign level2_sums[22:21] = pprod[5][12:11];


    // final add
    logic signed [23:0] add_result;
    assign add_result = level2_sums + {1'b0, level2_carries, 4'b0000};
    assign debug_output = add_result[21:0];
    assign overflow = add_result[21];
    assign result = add_result[20:8];      // Multiply result is the num_bits output bits plus two more: the R and S bits for rounding.
    assign round_loss = |add_result[7:0];

endmodule