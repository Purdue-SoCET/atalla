// lfc_ram_active_monitor.svh
`ifndef LFC_RAM_ACTIVE_MONITOR_SV
`define LFC_RAM_ACTIVE_MONITOR_SV

import uvm_pkg::*;
`include "uvm_macros.svh"
`include "lfc_if.sv"
`include "lfc_ram_transaction.sv"

// --- Replace these with your real types if needed ---
typedef virtual lfc_if lfc_ram_vif_t;
//typedef lfc_cpu_item       cpu_txn_t;

class lfc_ram_active_monitor extends uvm_monitor;
  `uvm_component_utils(lfc_ram_active_monitor)

  // analysis port to scoreboard/subscribers
  //uvm_analysis_port #(cpu_txn_t) ap;

  // optional: virtual interface handle
  lfc_cpu_vif_t vif;
  lfc_ram_transaction prev_tx;

  uvm_analysis_port#(lfc_ram_transaction) lfc_ap;

  function new(string name, uvm_component parent = null);
    super.new(name, parent);
    lfc_ap = new("lfc_ap", this);
  endfunction

  virtual function void build_phase(uvm_phase phase);
    super.build_phase(phase);
    //ap = new("ap", this);
    // optional: get VIF from config_db
    if(!uvm_config_db#(virtual lfc_if)::get(this, "", "lfc_vif", vif)) begin
      `uvm_fatal("Monitor", "No virtual interface specified for this monitor instance")
    end
  endfunction

  int has_run_once;
  virtual task run_phase(uvm_phase phase);
    super.run_phase(phase);
    prev_tx = lfc_ram_transaction::type_id::create("prev_tx");

    has_run_once = 0;
    forever begin
      lfc_ram_transaction tx;
      @(posedge vif.clk);
      tx = lfc_ram_transaction::type_id::create("tx");

      tx.ram_mem_data = vif.ram_mem_data;
      tx.ram_mem_complete = vif.ram_mem_complete;

      if(has_run_once > 0) begin // avoids an uninstantiated comparison
        if(tx.equal(prev.tx)) lfc_ap.write(tx);
      end

      prev_tx.copy(tx);
      if (has_run_once == 0) has_run_once++;
    end
  endtask

endclass

`endif // LFC_CPU_ACTIVE_MONITOR_SV
